/* 
Module to generate appropriate signals using the opcode and funct for R type instructions.
   1. RegDst - Which field of the instruction is the register to be written to
   2. RegWrite - Write to register file
   3. RegRead - Read from a register
   4. ALUSrc - The source for the second input to the ALU
   5. PCSrc - Source for PC (next instruction to be executed)
   6. MemRead - Read from the main memory
   7. MemWrite - Write to the main memory
   8. MemToReg - Source of write_data
   9. Branch -  When a branch/jump instruction is used
*/
module control_unit(
    output reg  RegRead,
                RegWrite,
                MemRead,
                MemWrite,
                RegDst, // 0: rt, 1: rd
                Branch,
                ALUSrc,
                PCSrc,
                MemToReg,
    input [5:0] opcode, funct
);

    always @(opcode, funct) 
    begin
	    // Reset all signals
        MemRead  = 1'b0;
        MemWrite = 1'b0;
        RegWrite = 1'b0;
        RegRead  = 1'b0;
        RegDst   = 1'b0;
        Branch   = 1'b0;
        ALUSrc   = 1'b0;
        PCSrc    = 1'b0;
        MemToReg = 1'b0;
		
        // R type
        if(opcode == 6'h0) begin
            RegDst = 1'b1;
            RegRead = 1'b1;
            // If NOT JR  - Jump Register
            if(funct != 6'h08) begin
                RegWrite = 1'b1;
            end
            // $display("RegWrite : %1b, RegDst : %1b, RegRead : %1b", RegWrite, RegDst, RegRead);
        end
        // LUI(load unsigned immediate) => no need to read any register => immediate value is written to a register
        else if(opcode == 6'b001111) begin
            RegWrite = 1'b1;
            ALUSrc   = 1'b1;
        end
        // If r-type, don't enter this block
        // For r-type, beq, bne, sb, sh and sw there is no need to register write
        else if(opcode != 6'h0 & opcode != 6'h4 & opcode != 6'h5 & opcode != 6'h28 & opcode != 6'h29 & opcode != 6'h2b) begin
            RegWrite = 1'b1;
        end
        // For branch instructions
        else if(opcode == 6'h4 | opcode == 6'h5) begin
            Branch   = 1'b1;
        end
        // For memory write operation
        // sb, sh and sw use memory to write
        else if(opcode != 6'h0 & (opcode == 6'h28 | opcode == 6'h29 | opcode == 6'h2b)) begin
            MemWrite = 1'b1;
            RegRead  = 1'b1;
            ALUSrc   = 1'b1;
        end
        // For memory read operation
        // lw, 
        else if(opcode != 6'h0 & (opcode == 6'h23))begin
            MemRead = 1'b1;
            ALUSrc  = 1'b1;
            MemToReg= 1'b1;
            RegRead = 1'b1;
        end
        // J type
        else
        begin
            PCSrc = 1'b1;
        end
    end
endmodule